reg q;
always @(posedge clk)
  q <= d;
