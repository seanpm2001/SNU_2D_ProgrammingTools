logic [1:0][2:0] my_pack[32];
