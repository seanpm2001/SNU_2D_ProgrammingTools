sequence S1;
    @(posedge clk) req ##1 gnt;
endsequence
