always_latch
    if (en) q <= d;
