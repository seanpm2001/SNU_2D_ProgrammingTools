always_comb begin
    tmp = b * b - 4 * a * c;
    no_root = (tmp < 0);
end

