always_ff @(posedge clk)
    count <= count + 1;
