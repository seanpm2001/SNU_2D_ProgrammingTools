-- Start of file
WRITE "CORRUPT" TO V://Root
IN FILE: hard.sys
X = 12
I = 1
FOR I in range(5)
	WRITE "TEST" TO "TEST"
WHILE X = X:
	WRITE "1" TO V://Root
begin buffer(6)
block []
block buffer
end block
end file
write "a" out
-- Just figuring out the syntax. Do not run this, as it won't work (100% guarantee) Virtual Hard Disk Language file.
-- File info:
-- Name: Test1
-- Extension: .VHDL (Virtual Hard Disk Language)
-- Language: VHDL (Virtual Hard Disk Language)
-- Stable? No
-- Functional? No
-- Version 1: September 8th 2019
-- Latest version: 1
-- End of file