logic [31:0] my_var;
